module mrd_ROM_fake (
	input clk,

	input [2:0]  factor,
	input [7:0]  wraddr,

	output logic signed [17:0] dout_real,
	output logic signed [17:0] dout_imag
);

// logic [59:0]  mem[0:255];
logic signed [29:0]  mem2_r[0:255];
logic signed [29:0]  mem2_i[0:255];
logic signed [29:0]  mem3_r[0:255];
logic signed [29:0]  mem3_i[0:255];
logic signed [29:0]  mem5_r[0:255];
logic signed [29:0]  mem5_i[0:255];
always@(posedge clk)
begin
	if (factor==3'd5)
	begin
		dout_real <= mem5_r[rdaddr];
		dout_imag <= mem5_i[rdaddr];
	end
	else if (factor==3'd3)
	begin
		dout_real <= mem3_r[rdaddr];
		dout_imag <= mem3_i[rdaddr];
	end
	else
	begin
		dout_real <= mem4_r[rdaddr];
		dout_imag <= mem4_i[rdaddr];
	end
end


assign mem4_r[0] = 18'd131072;
assign mem4_i[0] = 18'd0;
assign mem4_r[1] = 18'd131033;
assign mem4_i[1] = -18'd3217;
assign mem4_r[2] = 18'd130914;
assign mem4_i[2] = -18'd6431;
assign mem4_r[3] = 18'd130717;
assign mem4_i[3] = -18'd9642;
assign mem4_r[4] = 18'd130441;
assign mem4_i[4] = -18'd12847;
assign mem4_r[5] = 18'd130086;
assign mem4_i[5] = -18'd16045;
assign mem4_r[6] = 18'd129653;
assign mem4_i[6] = -18'd19232;
assign mem4_r[7] = 18'd129142;
assign mem4_i[7] = -18'd22408;
assign mem4_r[8] = 18'd128553;
assign mem4_i[8] = -18'd25571;
assign mem4_r[9] = 18'd127887;
assign mem4_i[9] = -18'd28718;
assign mem4_r[10] = 18'd127144;
assign mem4_i[10] = -18'd31848;
assign mem4_r[11] = 18'd126324;
assign mem4_i[11] = -18'd34959;
assign mem4_r[12] = 18'd125428;
assign mem4_i[12] = -18'd38048;
assign mem4_r[13] = 18'd124457;
assign mem4_i[13] = -18'd41115;
assign mem4_r[14] = 18'd123410;
assign mem4_i[14] = -18'd44157;
assign mem4_r[15] = 18'd122289;
assign mem4_i[15] = -18'd47172;
assign mem4_r[16] = 18'd121095;
assign mem4_i[16] = -18'd50159;
assign mem4_r[17] = 18'd119827;
assign mem4_i[17] = -18'd53116;
assign mem4_r[18] = 18'd118488;
assign mem4_i[18] = -18'd56041;
assign mem4_r[19] = 18'd117077;
assign mem4_i[19] = -18'd58931;
assign mem4_r[20] = 18'd115595;
assign mem4_i[20] = -18'd61787;
assign mem4_r[21] = 18'd114044;
assign mem4_i[21] = -18'd64605;
assign mem4_r[22] = 18'd112424;
assign mem4_i[22] = -18'd67384;
assign mem4_r[23] = 18'd110737;
assign mem4_i[23] = -18'd70123;
assign mem4_r[24] = 18'd108982;
assign mem4_i[24] = -18'd72820;
assign mem4_r[25] = 18'd107162;
assign mem4_i[25] = -18'd75472;
assign mem4_r[26] = 18'd105278;
assign mem4_i[26] = -18'd78079;
assign mem4_r[27] = 18'd103330;
assign mem4_i[27] = -18'd80640;
assign mem4_r[28] = 18'd101320;
assign mem4_i[28] = -18'd83151;
assign mem4_r[29] = 18'd99249;
assign mem4_i[29] = -18'd85613;
assign mem4_r[30] = 18'd97118;
assign mem4_i[30] = -18'd88023;
assign mem4_r[31] = 18'd94929;
assign mem4_i[31] = -18'd90379;
assign mem4_r[32] = 18'd92682;
assign mem4_i[32] = -18'd92682;
assign mem4_r[33] = 18'd90379;
assign mem4_i[33] = -18'd94929;
assign mem4_r[34] = 18'd88023;
assign mem4_i[34] = -18'd97118;
assign mem4_r[35] = 18'd85613;
assign mem4_i[35] = -18'd99249;
assign mem4_r[36] = 18'd83151;
assign mem4_i[36] = -18'd101320;
assign mem4_r[37] = 18'd80640;
assign mem4_i[37] = -18'd103330;
assign mem4_r[38] = 18'd78079;
assign mem4_i[38] = -18'd105278;
assign mem4_r[39] = 18'd75472;
assign mem4_i[39] = -18'd107162;
assign mem4_r[40] = 18'd72820;
assign mem4_i[40] = -18'd108982;
assign mem4_r[41] = 18'd70123;
assign mem4_i[41] = -18'd110737;
assign mem4_r[42] = 18'd67384;
assign mem4_i[42] = -18'd112424;
assign mem4_r[43] = 18'd64605;
assign mem4_i[43] = -18'd114044;
assign mem4_r[44] = 18'd61787;
assign mem4_i[44] = -18'd115595;
assign mem4_r[45] = 18'd58931;
assign mem4_i[45] = -18'd117077;
assign mem4_r[46] = 18'd56041;
assign mem4_i[46] = -18'd118488;
assign mem4_r[47] = 18'd53116;
assign mem4_i[47] = -18'd119827;
assign mem4_r[48] = 18'd50159;
assign mem4_i[48] = -18'd121095;
assign mem4_r[49] = 18'd47172;
assign mem4_i[49] = -18'd122289;
assign mem4_r[50] = 18'd44157;
assign mem4_i[50] = -18'd123410;
assign mem4_r[51] = 18'd41115;
assign mem4_i[51] = -18'd124457;
assign mem4_r[52] = 18'd38048;
assign mem4_i[52] = -18'd125428;
assign mem4_r[53] = 18'd34959;
assign mem4_i[53] = -18'd126324;
assign mem4_r[54] = 18'd31848;
assign mem4_i[54] = -18'd127144;
assign mem4_r[55] = 18'd28718;
assign mem4_i[55] = -18'd127887;
assign mem4_r[56] = 18'd25571;
assign mem4_i[56] = -18'd128553;
assign mem4_r[57] = 18'd22408;
assign mem4_i[57] = -18'd129142;
assign mem4_r[58] = 18'd19232;
assign mem4_i[58] = -18'd129653;
assign mem4_r[59] = 18'd16045;
assign mem4_i[59] = -18'd130086;
assign mem4_r[60] = 18'd12847;
assign mem4_i[60] = -18'd130441;
assign mem4_r[61] = 18'd9642;
assign mem4_i[61] = -18'd130717;
assign mem4_r[62] = 18'd6431;
assign mem4_i[62] = -18'd130914;
assign mem4_r[63] = 18'd3217;
assign mem4_i[63] = -18'd131033;
assign mem4_r[64] = 18'd0;
assign mem4_i[64] = -18'd131072;
assign mem4_r[65] = -18'd3217;
assign mem4_i[65] = -18'd131033;
assign mem4_r[66] = -18'd6431;
assign mem4_i[66] = -18'd130914;
assign mem4_r[67] = -18'd9642;
assign mem4_i[67] = -18'd130717;
assign mem4_r[68] = -18'd12847;
assign mem4_i[68] = -18'd130441;
assign mem4_r[69] = -18'd16045;
assign mem4_i[69] = -18'd130086;
assign mem4_r[70] = -18'd19232;
assign mem4_i[70] = -18'd129653;
assign mem4_r[71] = -18'd22408;
assign mem4_i[71] = -18'd129142;
assign mem4_r[72] = -18'd25571;
assign mem4_i[72] = -18'd128553;
assign mem4_r[73] = -18'd28718;
assign mem4_i[73] = -18'd127887;
assign mem4_r[74] = -18'd31848;
assign mem4_i[74] = -18'd127144;
assign mem4_r[75] = -18'd34959;
assign mem4_i[75] = -18'd126324;
assign mem4_r[76] = -18'd38048;
assign mem4_i[76] = -18'd125428;
assign mem4_r[77] = -18'd41115;
assign mem4_i[77] = -18'd124457;
assign mem4_r[78] = -18'd44157;
assign mem4_i[78] = -18'd123410;
assign mem4_r[79] = -18'd47172;
assign mem4_i[79] = -18'd122289;
assign mem4_r[80] = -18'd50159;
assign mem4_i[80] = -18'd121095;
assign mem4_r[81] = -18'd53116;
assign mem4_i[81] = -18'd119827;
assign mem4_r[82] = -18'd56041;
assign mem4_i[82] = -18'd118488;
assign mem4_r[83] = -18'd58931;
assign mem4_i[83] = -18'd117077;
assign mem4_r[84] = -18'd61787;
assign mem4_i[84] = -18'd115595;
assign mem4_r[85] = -18'd64605;
assign mem4_i[85] = -18'd114044;
assign mem4_r[86] = -18'd67384;
assign mem4_i[86] = -18'd112424;
assign mem4_r[87] = -18'd70123;
assign mem4_i[87] = -18'd110737;
assign mem4_r[88] = -18'd72820;
assign mem4_i[88] = -18'd108982;
assign mem4_r[89] = -18'd75472;
assign mem4_i[89] = -18'd107162;
assign mem4_r[90] = -18'd78079;
assign mem4_i[90] = -18'd105278;
assign mem4_r[91] = -18'd80640;
assign mem4_i[91] = -18'd103330;
assign mem4_r[92] = -18'd83151;
assign mem4_i[92] = -18'd101320;
assign mem4_r[93] = -18'd85613;
assign mem4_i[93] = -18'd99249;
assign mem4_r[94] = -18'd88023;
assign mem4_i[94] = -18'd97118;
assign mem4_r[95] = -18'd90379;
assign mem4_i[95] = -18'd94929;
assign mem4_r[96] = -18'd92682;
assign mem4_i[96] = -18'd92682;
assign mem4_r[97] = -18'd94929;
assign mem4_i[97] = -18'd90379;
assign mem4_r[98] = -18'd97118;
assign mem4_i[98] = -18'd88023;
assign mem4_r[99] = -18'd99249;
assign mem4_i[99] = -18'd85613;
assign mem4_r[100] = -18'd101320;
assign mem4_i[100] = -18'd83151;
assign mem4_r[101] = -18'd103330;
assign mem4_i[101] = -18'd80640;
assign mem4_r[102] = -18'd105278;
assign mem4_i[102] = -18'd78079;
assign mem4_r[103] = -18'd107162;
assign mem4_i[103] = -18'd75472;
assign mem4_r[104] = -18'd108982;
assign mem4_i[104] = -18'd72820;
assign mem4_r[105] = -18'd110737;
assign mem4_i[105] = -18'd70123;
assign mem4_r[106] = -18'd112424;
assign mem4_i[106] = -18'd67384;
assign mem4_r[107] = -18'd114044;
assign mem4_i[107] = -18'd64605;
assign mem4_r[108] = -18'd115595;
assign mem4_i[108] = -18'd61787;
assign mem4_r[109] = -18'd117077;
assign mem4_i[109] = -18'd58931;
assign mem4_r[110] = -18'd118488;
assign mem4_i[110] = -18'd56041;
assign mem4_r[111] = -18'd119827;
assign mem4_i[111] = -18'd53116;
assign mem4_r[112] = -18'd121095;
assign mem4_i[112] = -18'd50159;
assign mem4_r[113] = -18'd122289;
assign mem4_i[113] = -18'd47172;
assign mem4_r[114] = -18'd123410;
assign mem4_i[114] = -18'd44157;
assign mem4_r[115] = -18'd124457;
assign mem4_i[115] = -18'd41115;
assign mem4_r[116] = -18'd125428;
assign mem4_i[116] = -18'd38048;
assign mem4_r[117] = -18'd126324;
assign mem4_i[117] = -18'd34959;
assign mem4_r[118] = -18'd127144;
assign mem4_i[118] = -18'd31848;
assign mem4_r[119] = -18'd127887;
assign mem4_i[119] = -18'd28718;
assign mem4_r[120] = -18'd128553;
assign mem4_i[120] = -18'd25571;
assign mem4_r[121] = -18'd129142;
assign mem4_i[121] = -18'd22408;
assign mem4_r[122] = -18'd129653;
assign mem4_i[122] = -18'd19232;
assign mem4_r[123] = -18'd130086;
assign mem4_i[123] = -18'd16045;
assign mem4_r[124] = -18'd130441;
assign mem4_i[124] = -18'd12847;
assign mem4_r[125] = -18'd130717;
assign mem4_i[125] = -18'd9642;
assign mem4_r[126] = -18'd130914;
assign mem4_i[126] = -18'd6431;
assign mem4_r[127] = -18'd131033;
assign mem4_i[127] = -18'd3217;
assign mem4_r[128] = -18'd131072;
assign mem4_i[128] = 18'd0;
assign mem4_r[129] = -18'd131033;
assign mem4_i[129] = 18'd3217;
assign mem4_r[130] = -18'd130914;
assign mem4_i[130] = 18'd6431;
assign mem4_r[131] = -18'd130717;
assign mem4_i[131] = 18'd9642;
assign mem4_r[132] = -18'd130441;
assign mem4_i[132] = 18'd12847;
assign mem4_r[133] = -18'd130086;
assign mem4_i[133] = 18'd16045;
assign mem4_r[134] = -18'd129653;
assign mem4_i[134] = 18'd19232;
assign mem4_r[135] = -18'd129142;
assign mem4_i[135] = 18'd22408;
assign mem4_r[136] = -18'd128553;
assign mem4_i[136] = 18'd25571;
assign mem4_r[137] = -18'd127887;
assign mem4_i[137] = 18'd28718;
assign mem4_r[138] = -18'd127144;
assign mem4_i[138] = 18'd31848;
assign mem4_r[139] = -18'd126324;
assign mem4_i[139] = 18'd34959;
assign mem4_r[140] = -18'd125428;
assign mem4_i[140] = 18'd38048;
assign mem4_r[141] = -18'd124457;
assign mem4_i[141] = 18'd41115;
assign mem4_r[142] = -18'd123410;
assign mem4_i[142] = 18'd44157;
assign mem4_r[143] = -18'd122289;
assign mem4_i[143] = 18'd47172;
assign mem4_r[144] = -18'd121095;
assign mem4_i[144] = 18'd50159;
assign mem4_r[145] = -18'd119827;
assign mem4_i[145] = 18'd53116;
assign mem4_r[146] = -18'd118488;
assign mem4_i[146] = 18'd56041;
assign mem4_r[147] = -18'd117077;
assign mem4_i[147] = 18'd58931;
assign mem4_r[148] = -18'd115595;
assign mem4_i[148] = 18'd61787;
assign mem4_r[149] = -18'd114044;
assign mem4_i[149] = 18'd64605;
assign mem4_r[150] = -18'd112424;
assign mem4_i[150] = 18'd67384;
assign mem4_r[151] = -18'd110737;
assign mem4_i[151] = 18'd70123;
assign mem4_r[152] = -18'd108982;
assign mem4_i[152] = 18'd72820;
assign mem4_r[153] = -18'd107162;
assign mem4_i[153] = 18'd75472;
assign mem4_r[154] = -18'd105278;
assign mem4_i[154] = 18'd78079;
assign mem4_r[155] = -18'd103330;
assign mem4_i[155] = 18'd80640;
assign mem4_r[156] = -18'd101320;
assign mem4_i[156] = 18'd83151;
assign mem4_r[157] = -18'd99249;
assign mem4_i[157] = 18'd85613;
assign mem4_r[158] = -18'd97118;
assign mem4_i[158] = 18'd88023;
assign mem4_r[159] = -18'd94929;
assign mem4_i[159] = 18'd90379;
assign mem4_r[160] = -18'd92682;
assign mem4_i[160] = 18'd92682;
assign mem4_r[161] = -18'd90379;
assign mem4_i[161] = 18'd94929;
assign mem4_r[162] = -18'd88023;
assign mem4_i[162] = 18'd97118;
assign mem4_r[163] = -18'd85613;
assign mem4_i[163] = 18'd99249;
assign mem4_r[164] = -18'd83151;
assign mem4_i[164] = 18'd101320;
assign mem4_r[165] = -18'd80640;
assign mem4_i[165] = 18'd103330;
assign mem4_r[166] = -18'd78079;
assign mem4_i[166] = 18'd105278;
assign mem4_r[167] = -18'd75472;
assign mem4_i[167] = 18'd107162;
assign mem4_r[168] = -18'd72820;
assign mem4_i[168] = 18'd108982;
assign mem4_r[169] = -18'd70123;
assign mem4_i[169] = 18'd110737;
assign mem4_r[170] = -18'd67384;
assign mem4_i[170] = 18'd112424;
assign mem4_r[171] = -18'd64605;
assign mem4_i[171] = 18'd114044;
assign mem4_r[172] = -18'd61787;
assign mem4_i[172] = 18'd115595;
assign mem4_r[173] = -18'd58931;
assign mem4_i[173] = 18'd117077;
assign mem4_r[174] = -18'd56041;
assign mem4_i[174] = 18'd118488;
assign mem4_r[175] = -18'd53116;
assign mem4_i[175] = 18'd119827;
assign mem4_r[176] = -18'd50159;
assign mem4_i[176] = 18'd121095;
assign mem4_r[177] = -18'd47172;
assign mem4_i[177] = 18'd122289;
assign mem4_r[178] = -18'd44157;
assign mem4_i[178] = 18'd123410;
assign mem4_r[179] = -18'd41115;
assign mem4_i[179] = 18'd124457;
assign mem4_r[180] = -18'd38048;
assign mem4_i[180] = 18'd125428;
assign mem4_r[181] = -18'd34959;
assign mem4_i[181] = 18'd126324;
assign mem4_r[182] = -18'd31848;
assign mem4_i[182] = 18'd127144;
assign mem4_r[183] = -18'd28718;
assign mem4_i[183] = 18'd127887;
assign mem4_r[184] = -18'd25571;
assign mem4_i[184] = 18'd128553;
assign mem4_r[185] = -18'd22408;
assign mem4_i[185] = 18'd129142;
assign mem4_r[186] = -18'd19232;
assign mem4_i[186] = 18'd129653;
assign mem4_r[187] = -18'd16045;
assign mem4_i[187] = 18'd130086;
assign mem4_r[188] = -18'd12847;
assign mem4_i[188] = 18'd130441;
assign mem4_r[189] = -18'd9642;
assign mem4_i[189] = 18'd130717;
assign mem4_r[190] = -18'd6431;
assign mem4_i[190] = 18'd130914;
assign mem4_r[191] = -18'd3217;
assign mem4_i[191] = 18'd131033;
assign mem4_r[192] = 18'd0;
assign mem4_i[192] = 18'd131072;
assign mem4_r[193] = 18'd3217;
assign mem4_i[193] = 18'd131033;
assign mem4_r[194] = 18'd6431;
assign mem4_i[194] = 18'd130914;
assign mem4_r[195] = 18'd9642;
assign mem4_i[195] = 18'd130717;
assign mem4_r[196] = 18'd12847;
assign mem4_i[196] = 18'd130441;
assign mem4_r[197] = 18'd16045;
assign mem4_i[197] = 18'd130086;
assign mem4_r[198] = 18'd19232;
assign mem4_i[198] = 18'd129653;
assign mem4_r[199] = 18'd22408;
assign mem4_i[199] = 18'd129142;
assign mem4_r[200] = 18'd25571;
assign mem4_i[200] = 18'd128553;
assign mem4_r[201] = 18'd28718;
assign mem4_i[201] = 18'd127887;
assign mem4_r[202] = 18'd31848;
assign mem4_i[202] = 18'd127144;
assign mem4_r[203] = 18'd34959;
assign mem4_i[203] = 18'd126324;
assign mem4_r[204] = 18'd38048;
assign mem4_i[204] = 18'd125428;
assign mem4_r[205] = 18'd41115;
assign mem4_i[205] = 18'd124457;
assign mem4_r[206] = 18'd44157;
assign mem4_i[206] = 18'd123410;
assign mem4_r[207] = 18'd47172;
assign mem4_i[207] = 18'd122289;
assign mem4_r[208] = 18'd50159;
assign mem4_i[208] = 18'd121095;
assign mem4_r[209] = 18'd53116;
assign mem4_i[209] = 18'd119827;
assign mem4_r[210] = 18'd56041;
assign mem4_i[210] = 18'd118488;
assign mem4_r[211] = 18'd58931;
assign mem4_i[211] = 18'd117077;
assign mem4_r[212] = 18'd61787;
assign mem4_i[212] = 18'd115595;
assign mem4_r[213] = 18'd64605;
assign mem4_i[213] = 18'd114044;
assign mem4_r[214] = 18'd67384;
assign mem4_i[214] = 18'd112424;
assign mem4_r[215] = 18'd70123;
assign mem4_i[215] = 18'd110737;
assign mem4_r[216] = 18'd72820;
assign mem4_i[216] = 18'd108982;
assign mem4_r[217] = 18'd75472;
assign mem4_i[217] = 18'd107162;
assign mem4_r[218] = 18'd78079;
assign mem4_i[218] = 18'd105278;
assign mem4_r[219] = 18'd80640;
assign mem4_i[219] = 18'd103330;
assign mem4_r[220] = 18'd83151;
assign mem4_i[220] = 18'd101320;
assign mem4_r[221] = 18'd85613;
assign mem4_i[221] = 18'd99249;
assign mem4_r[222] = 18'd88023;
assign mem4_i[222] = 18'd97118;
assign mem4_r[223] = 18'd90379;
assign mem4_i[223] = 18'd94929;
assign mem4_r[224] = 18'd92682;
assign mem4_i[224] = 18'd92682;
assign mem4_r[225] = 18'd94929;
assign mem4_i[225] = 18'd90379;
assign mem4_r[226] = 18'd97118;
assign mem4_i[226] = 18'd88023;
assign mem4_r[227] = 18'd99249;
assign mem4_i[227] = 18'd85613;
assign mem4_r[228] = 18'd101320;
assign mem4_i[228] = 18'd83151;
assign mem4_r[229] = 18'd103330;
assign mem4_i[229] = 18'd80640;
assign mem4_r[230] = 18'd105278;
assign mem4_i[230] = 18'd78079;
assign mem4_r[231] = 18'd107162;
assign mem4_i[231] = 18'd75472;
assign mem4_r[232] = 18'd108982;
assign mem4_i[232] = 18'd72820;
assign mem4_r[233] = 18'd110737;
assign mem4_i[233] = 18'd70123;
assign mem4_r[234] = 18'd112424;
assign mem4_i[234] = 18'd67384;
assign mem4_r[235] = 18'd114044;
assign mem4_i[235] = 18'd64605;
assign mem4_r[236] = 18'd115595;
assign mem4_i[236] = 18'd61787;
assign mem4_r[237] = 18'd117077;
assign mem4_i[237] = 18'd58931;
assign mem4_r[238] = 18'd118488;
assign mem4_i[238] = 18'd56041;
assign mem4_r[239] = 18'd119827;
assign mem4_i[239] = 18'd53116;
assign mem4_r[240] = 18'd121095;
assign mem4_i[240] = 18'd50159;
assign mem4_r[241] = 18'd122289;
assign mem4_i[241] = 18'd47172;
assign mem4_r[242] = 18'd123410;
assign mem4_i[242] = 18'd44157;
assign mem4_r[243] = 18'd124457;
assign mem4_i[243] = 18'd41115;
assign mem4_r[244] = 18'd125428;
assign mem4_i[244] = 18'd38048;
assign mem4_r[245] = 18'd126324;
assign mem4_i[245] = 18'd34959;
assign mem4_r[246] = 18'd127144;
assign mem4_i[246] = 18'd31848;
assign mem4_r[247] = 18'd127887;
assign mem4_i[247] = 18'd28718;
assign mem4_r[248] = 18'd128553;
assign mem4_i[248] = 18'd25571;
assign mem4_r[249] = 18'd129142;
assign mem4_i[249] = 18'd22408;
assign mem4_r[250] = 18'd129653;
assign mem4_i[250] = 18'd19232;
assign mem4_r[251] = 18'd130086;
assign mem4_i[251] = 18'd16045;
assign mem4_r[252] = 18'd130441;
assign mem4_i[252] = 18'd12847;
assign mem4_r[253] = 18'd130717;
assign mem4_i[253] = 18'd9642;
assign mem4_r[254] = 18'd130914;
assign mem4_i[254] = 18'd6431;
assign mem4_r[255] = 18'd131033;
assign mem4_i[255] = 18'd3217;




endmodule