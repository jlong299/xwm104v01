
module lpm_mult_18_mrd (
	dataa,
	datab,
	clock,
	result);	

	input	[17:0]	dataa;
	input	[17:0]	datab;
	input		clock;
	output	[35:0]	result;
endmodule
