
module lpm_mult_16_mrd (
	dataa,
	datab,
	clock,
	result);	

	input	[15:0]	dataa;
	input	[15:0]	datab;
	input		clock;
	output	[31:0]	result;
endmodule
