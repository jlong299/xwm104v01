
module mrd_ROM_Init (
	address,
	clock,
	q);	

	input	[6:0]	address;
	input		clock;
	output	[63:0]	q;
endmodule
