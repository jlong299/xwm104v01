
module lpm_mult_1816_mrd (
	dataa,
	datab,
	clock,
	result);	

	input	[17:0]	dataa;
	input	[15:0]	datab;
	input		clock;
	output	[33:0]	result;
endmodule
