module mrd_ROM_fake (
	input clk,

	input [2:0]  factor,
	input [7:0]  rdaddr,

	output logic signed [17:0] dout_real,
	output logic signed [17:0] dout_imag
);

// logic [59:0]  mem[0:255];
logic signed [29:0]  mem2_r[0:255];
logic signed [29:0]  mem2_i[0:255];
logic signed [29:0]  mem3_r[0:255];
logic signed [29:0]  mem3_i[0:255];
logic signed [29:0]  mem5_r[0:255];
logic signed [29:0]  mem5_i[0:255];
always@(posedge clk)
begin
	if (factor==3'd5)
	begin
		dout_real <= mem5_r[rdaddr];
		dout_imag <= mem5_i[rdaddr];
	end
	else if (factor==3'd3)
	begin
		dout_real <= mem3_r[rdaddr];
		dout_imag <= mem3_i[rdaddr];
	end
	else
	begin
		dout_real <= mem2_r[rdaddr];
		dout_imag <= mem2_i[rdaddr];
	end
end


assign mem5_r[0] = 18'd65536;
assign mem5_i[0] = 18'd0;
assign mem5_r[1] = 18'd63477;
assign mem5_i[1] = -18'd16298;
assign mem5_r[2] = 18'd57430;
assign mem5_i[2] = -18'd31572;
assign mem5_r[3] = 18'd47774;
assign mem5_i[3] = -18'd44862;
assign mem5_r[4] = 18'd35116;
assign mem5_i[4] = -18'd55334;
assign mem5_r[5] = 18'd20252;
assign mem5_i[5] = -18'd62328;
assign mem5_r[6] = 18'd4115;
assign mem5_i[6] = -18'd65407;
assign mem5_r[7] = -18'd12280;
assign mem5_i[7] = -18'd64375;
assign mem5_r[8] = -18'd27904;
assign mem5_i[8] = -18'd59299;
assign mem5_r[9] = -18'd41774;
assign mem5_i[9] = -18'd50496;
assign mem5_r[10] = -18'd53020;
assign mem5_i[10] = -18'd38521;
assign mem5_r[11] = -18'd60934;
assign mem5_i[11] = -18'd24125;
assign mem5_r[12] = -18'd65019;
assign mem5_i[12] = -18'd8214;
assign mem5_r[13] = -18'd65019;
assign mem5_i[13] = 18'd8214;
assign mem5_r[14] = -18'd60934;
assign mem5_i[14] = 18'd24125;
assign mem5_r[15] = -18'd53020;
assign mem5_i[15] = 18'd38521;
assign mem5_r[16] = -18'd41774;
assign mem5_i[16] = 18'd50496;
assign mem5_r[17] = -18'd27904;
assign mem5_i[17] = 18'd59299;
assign mem5_r[18] = -18'd12280;
assign mem5_i[18] = 18'd64375;
assign mem5_r[19] = 18'd4115;
assign mem5_i[19] = 18'd65407;
assign mem5_r[20] = 18'd20252;
assign mem5_i[20] = 18'd62328;
assign mem5_r[21] = 18'd35116;
assign mem5_i[21] = 18'd55334;
assign mem5_r[22] = 18'd47774;
assign mem5_i[22] = 18'd44862;
assign mem5_r[23] = 18'd57430;
assign mem5_i[23] = 18'd31572;
assign mem5_r[24] = 18'd63477;
assign mem5_i[24] = 18'd16298;


assign mem3_r[0] = 18'd65536;
assign mem3_i[0] = 18'd0;
assign mem3_r[1] = 18'd65514;
assign mem3_i[1] = -18'd1694;
assign mem3_r[2] = 18'd65448;
assign mem3_i[2] = -18'd3388;
assign mem3_r[3] = 18'd65339;
assign mem3_i[3] = -18'd5079;
assign mem3_r[4] = 18'd65186;
assign mem3_i[4] = -18'd6766;
assign mem3_r[5] = 18'd64989;
assign mem3_i[5] = -18'd8449;
assign mem3_r[6] = 18'd64749;
assign mem3_i[6] = -18'd10127;
assign mem3_r[7] = 18'd64465;
assign mem3_i[7] = -18'd11797;
assign mem3_r[8] = 18'd64139;
assign mem3_i[8] = -18'd13460;
assign mem3_r[9] = 18'd63769;
assign mem3_i[9] = -18'd15114;
assign mem3_r[10] = 18'd63357;
assign mem3_i[10] = -18'd16757;
assign mem3_r[11] = 18'd62903;
assign mem3_i[11] = -18'd18390;
assign mem3_r[12] = 18'd62407;
assign mem3_i[12] = -18'd20010;
assign mem3_r[13] = 18'd61868;
assign mem3_i[13] = -18'd21617;
assign mem3_r[14] = 18'd61289;
assign mem3_i[14] = -18'd23209;
assign mem3_r[15] = 18'd60668;
assign mem3_i[15] = -18'd24786;
assign mem3_r[16] = 18'd60007;
assign mem3_i[16] = -18'd26346;
assign mem3_r[17] = 18'd59306;
assign mem3_i[17] = -18'd27889;
assign mem3_r[18] = 18'd58565;
assign mem3_i[18] = -18'd29413;
assign mem3_r[19] = 18'd57785;
assign mem3_i[19] = -18'd30917;
assign mem3_r[20] = 18'd56966;
assign mem3_i[20] = -18'd32400;
assign mem3_r[21] = 18'd56110;
assign mem3_i[21] = -18'd33862;
assign mem3_r[22] = 18'd55216;
assign mem3_i[22] = -18'd35302;
assign mem3_r[23] = 18'd54284;
assign mem3_i[23] = -18'd36717;
assign mem3_r[24] = 18'd53317;
assign mem3_i[24] = -18'd38109;
assign mem3_r[25] = 18'd52314;
assign mem3_i[25] = -18'd39474;
assign mem3_r[26] = 18'd51276;
assign mem3_i[26] = -18'd40814;
assign mem3_r[27] = 18'd50203;
assign mem3_i[27] = -18'd42126;
assign mem3_r[28] = 18'd49098;
assign mem3_i[28] = -18'd43410;
assign mem3_r[29] = 18'd47959;
assign mem3_i[29] = -18'd44664;
assign mem3_r[30] = 18'd46788;
assign mem3_i[30] = -18'd45889;
assign mem3_r[31] = 18'd45586;
assign mem3_i[31] = -18'd47084;
assign mem3_r[32] = 18'd44354;
assign mem3_i[32] = -18'd48247;
assign mem3_r[33] = 18'd43091;
assign mem3_i[33] = -18'd49377;
assign mem3_r[34] = 18'd41800;
assign mem3_i[34] = -18'd50475;
assign mem3_r[35] = 18'd40481;
assign mem3_i[35] = -18'd51539;
assign mem3_r[36] = 18'd39135;
assign mem3_i[36] = -18'd52568;
assign mem3_r[37] = 18'd37763;
assign mem3_i[37] = -18'd53562;
assign mem3_r[38] = 18'd36366;
assign mem3_i[38] = -18'd54521;
assign mem3_r[39] = 18'd34944;
assign mem3_i[39] = -18'd55443;
assign mem3_r[40] = 18'd33499;
assign mem3_i[40] = -18'd56327;
assign mem3_r[41] = 18'd32032;
assign mem3_i[41] = -18'd57175;
assign mem3_r[42] = 18'd30543;
assign mem3_i[42] = -18'd57984;
assign mem3_r[43] = 18'd29033;
assign mem3_i[43] = -18'd58754;
assign mem3_r[44] = 18'd27505;
assign mem3_i[44] = -18'd59485;
assign mem3_r[45] = 18'd25957;
assign mem3_i[45] = -18'd60176;
assign mem3_r[46] = 18'd24393;
assign mem3_i[46] = -18'd60827;
assign mem3_r[47] = 18'd22812;
assign mem3_i[47] = -18'd61438;
assign mem3_r[48] = 18'd21216;
assign mem3_i[48] = -18'd62007;
assign mem3_r[49] = 18'd19606;
assign mem3_i[49] = -18'd62535;
assign mem3_r[50] = 18'd17983;
assign mem3_i[50] = -18'd63021;
assign mem3_r[51] = 18'd16347;
assign mem3_i[51] = -18'd63464;
assign mem3_r[52] = 18'd14701;
assign mem3_i[52] = -18'd63866;
assign mem3_r[53] = 18'd13045;
assign mem3_i[53] = -18'd64225;
assign mem3_r[54] = 18'd11380;
assign mem3_i[54] = -18'd64540;
assign mem3_r[55] = 18'd9708;
assign mem3_i[55] = -18'd64813;
assign mem3_r[56] = 18'd8029;
assign mem3_i[56] = -18'd65042;
assign mem3_r[57] = 18'd6345;
assign mem3_i[57] = -18'd65228;
assign mem3_r[58] = 18'd4656;
assign mem3_i[58] = -18'd65370;
assign mem3_r[59] = 18'd2964;
assign mem3_i[59] = -18'd65469;
assign mem3_r[60] = 18'd1271;
assign mem3_i[60] = -18'd65524;
assign mem3_r[61] = -18'd424;
assign mem3_i[61] = -18'd65535;
assign mem3_r[62] = -18'd2118;
assign mem3_i[62] = -18'd65502;
assign mem3_r[63] = -18'd3811;
assign mem3_i[63] = -18'd65425;
assign mem3_r[64] = -18'd5501;
assign mem3_i[64] = -18'd65305;
assign mem3_r[65] = -18'd7187;
assign mem3_i[65] = -18'd65141;
assign mem3_r[66] = -18'd8869;
assign mem3_i[66] = -18'd64933;
assign mem3_r[67] = -18'd10545;
assign mem3_i[67] = -18'd64682;
assign mem3_r[68] = -18'd12214;
assign mem3_i[68] = -18'd64388;
assign mem3_r[69] = -18'd13874;
assign mem3_i[69] = -18'd64051;
assign mem3_r[70] = -18'd15526;
assign mem3_i[70] = -18'd63670;
assign mem3_r[71] = -18'd17166;
assign mem3_i[71] = -18'd63248;
assign mem3_r[72] = -18'd18796;
assign mem3_i[72] = -18'd62783;
assign mem3_r[73] = -18'd20413;
assign mem3_i[73] = -18'd62276;
assign mem3_r[74] = -18'd22016;
assign mem3_i[74] = -18'd61727;
assign mem3_r[75] = -18'd23605;
assign mem3_i[75] = -18'd61137;
assign mem3_r[76] = -18'd25177;
assign mem3_i[76] = -18'd60507;
assign mem3_r[77] = -18'd26733;
assign mem3_i[77] = -18'd59836;
assign mem3_r[78] = -18'd28271;
assign mem3_i[78] = -18'd59124;
assign mem3_r[79] = -18'd29790;
assign mem3_i[79] = -18'd58374;
assign mem3_r[80] = -18'd31290;
assign mem3_i[80] = -18'd57584;
assign mem3_r[81] = -18'd32768;
assign mem3_i[81] = -18'd56756;
assign mem3_r[82] = -18'd34224;
assign mem3_i[82] = -18'd55890;
assign mem3_r[83] = -18'd35658;
assign mem3_i[83] = -18'd54986;
assign mem3_r[84] = -18'd37068;
assign mem3_i[84] = -18'd54046;
assign mem3_r[85] = -18'd38453;
assign mem3_i[85] = -18'd53069;
assign mem3_r[86] = -18'd39812;
assign mem3_i[86] = -18'd52058;
assign mem3_r[87] = -18'd41144;
assign mem3_i[87] = -18'd51011;
assign mem3_r[88] = -18'd42449;
assign mem3_i[88] = -18'd49930;
assign mem3_r[89] = -18'd43726;
assign mem3_i[89] = -18'd48816;
assign mem3_r[90] = -18'd44974;
assign mem3_i[90] = -18'd47669;
assign mem3_r[91] = -18'd46191;
assign mem3_i[91] = -18'd46490;
assign mem3_r[92] = -18'd47377;
assign mem3_i[92] = -18'd45281;
assign mem3_r[93] = -18'd48532;
assign mem3_i[93] = -18'd44041;
assign mem3_r[94] = -18'd49655;
assign mem3_i[94] = -18'd42771;
assign mem3_r[95] = -18'd50744;
assign mem3_i[95] = -18'd41473;
assign mem3_r[96] = -18'd51799;
assign mem3_i[96] = -18'd40147;
assign mem3_r[97] = -18'd52820;
assign mem3_i[97] = -18'd38795;
assign mem3_r[98] = -18'd53805;
assign mem3_i[98] = -18'd37416;
assign mem3_r[99] = -18'd54755;
assign mem3_i[99] = -18'd36013;
assign mem3_r[100] = -18'd55667;
assign mem3_i[100] = -18'd34585;
assign mem3_r[101] = -18'd56543;
assign mem3_i[101] = -18'd33134;
assign mem3_r[102] = -18'd57381;
assign mem3_i[102] = -18'd31661;
assign mem3_r[103] = -18'd58180;
assign mem3_i[103] = -18'd30167;
assign mem3_r[104] = -18'd58940;
assign mem3_i[104] = -18'd28653;
assign mem3_r[105] = -18'd59662;
assign mem3_i[105] = -18'd27119;
assign mem3_r[106] = -18'd60343;
assign mem3_i[106] = -18'd25568;
assign mem3_r[107] = -18'd60984;
assign mem3_i[107] = -18'd23999;
assign mem3_r[108] = -18'd61584;
assign mem3_i[108] = -18'd22415;
assign mem3_r[109] = -18'd62143;
assign mem3_i[109] = -18'd20815;
assign mem3_r[110] = -18'd62660;
assign mem3_i[110] = -18'd19201;
assign mem3_r[111] = -18'd63135;
assign mem3_i[111] = -18'd17575;
assign mem3_r[112] = -18'd63569;
assign mem3_i[112] = -18'd15937;
assign mem3_r[113] = -18'd63960;
assign mem3_i[113] = -18'd14288;
assign mem3_r[114] = -18'd64308;
assign mem3_i[114] = -18'd12630;
assign mem3_r[115] = -18'd64613;
assign mem3_i[115] = -18'd10963;
assign mem3_r[116] = -18'd64874;
assign mem3_i[116] = -18'd9289;
assign mem3_r[117] = -18'd65093;
assign mem3_i[117] = -18'd7608;
assign mem3_r[118] = -18'd65268;
assign mem3_i[118] = -18'd5923;
assign mem3_r[119] = -18'd65399;
assign mem3_i[119] = -18'd4233;
assign mem3_r[120] = -18'd65487;
assign mem3_i[120] = -18'd2541;
assign mem3_r[121] = -18'd65531;
assign mem3_i[121] = -18'd847;
assign mem3_r[122] = -18'd65531;
assign mem3_i[122] = 18'd847;
assign mem3_r[123] = -18'd65487;
assign mem3_i[123] = 18'd2541;
assign mem3_r[124] = -18'd65399;
assign mem3_i[124] = 18'd4233;
assign mem3_r[125] = -18'd65268;
assign mem3_i[125] = 18'd5923;
assign mem3_r[126] = -18'd65093;
assign mem3_i[126] = 18'd7608;
assign mem3_r[127] = -18'd64874;
assign mem3_i[127] = 18'd9289;
assign mem3_r[128] = -18'd64613;
assign mem3_i[128] = 18'd10963;
assign mem3_r[129] = -18'd64308;
assign mem3_i[129] = 18'd12630;
assign mem3_r[130] = -18'd63960;
assign mem3_i[130] = 18'd14288;
assign mem3_r[131] = -18'd63569;
assign mem3_i[131] = 18'd15937;
assign mem3_r[132] = -18'd63135;
assign mem3_i[132] = 18'd17575;
assign mem3_r[133] = -18'd62660;
assign mem3_i[133] = 18'd19201;
assign mem3_r[134] = -18'd62143;
assign mem3_i[134] = 18'd20815;
assign mem3_r[135] = -18'd61584;
assign mem3_i[135] = 18'd22415;
assign mem3_r[136] = -18'd60984;
assign mem3_i[136] = 18'd23999;
assign mem3_r[137] = -18'd60343;
assign mem3_i[137] = 18'd25568;
assign mem3_r[138] = -18'd59662;
assign mem3_i[138] = 18'd27119;
assign mem3_r[139] = -18'd58940;
assign mem3_i[139] = 18'd28653;
assign mem3_r[140] = -18'd58180;
assign mem3_i[140] = 18'd30167;
assign mem3_r[141] = -18'd57381;
assign mem3_i[141] = 18'd31661;
assign mem3_r[142] = -18'd56543;
assign mem3_i[142] = 18'd33134;
assign mem3_r[143] = -18'd55667;
assign mem3_i[143] = 18'd34585;
assign mem3_r[144] = -18'd54755;
assign mem3_i[144] = 18'd36013;
assign mem3_r[145] = -18'd53805;
assign mem3_i[145] = 18'd37416;
assign mem3_r[146] = -18'd52820;
assign mem3_i[146] = 18'd38795;
assign mem3_r[147] = -18'd51799;
assign mem3_i[147] = 18'd40147;
assign mem3_r[148] = -18'd50744;
assign mem3_i[148] = 18'd41473;
assign mem3_r[149] = -18'd49655;
assign mem3_i[149] = 18'd42771;
assign mem3_r[150] = -18'd48532;
assign mem3_i[150] = 18'd44041;
assign mem3_r[151] = -18'd47377;
assign mem3_i[151] = 18'd45281;
assign mem3_r[152] = -18'd46191;
assign mem3_i[152] = 18'd46490;
assign mem3_r[153] = -18'd44974;
assign mem3_i[153] = 18'd47669;
assign mem3_r[154] = -18'd43726;
assign mem3_i[154] = 18'd48816;
assign mem3_r[155] = -18'd42449;
assign mem3_i[155] = 18'd49930;
assign mem3_r[156] = -18'd41144;
assign mem3_i[156] = 18'd51011;
assign mem3_r[157] = -18'd39812;
assign mem3_i[157] = 18'd52058;
assign mem3_r[158] = -18'd38453;
assign mem3_i[158] = 18'd53069;
assign mem3_r[159] = -18'd37068;
assign mem3_i[159] = 18'd54046;
assign mem3_r[160] = -18'd35658;
assign mem3_i[160] = 18'd54986;
assign mem3_r[161] = -18'd34224;
assign mem3_i[161] = 18'd55890;
assign mem3_r[162] = -18'd32768;
assign mem3_i[162] = 18'd56756;
assign mem3_r[163] = -18'd31290;
assign mem3_i[163] = 18'd57584;
assign mem3_r[164] = -18'd29790;
assign mem3_i[164] = 18'd58374;
assign mem3_r[165] = -18'd28271;
assign mem3_i[165] = 18'd59124;
assign mem3_r[166] = -18'd26733;
assign mem3_i[166] = 18'd59836;
assign mem3_r[167] = -18'd25177;
assign mem3_i[167] = 18'd60507;
assign mem3_r[168] = -18'd23605;
assign mem3_i[168] = 18'd61137;
assign mem3_r[169] = -18'd22016;
assign mem3_i[169] = 18'd61727;
assign mem3_r[170] = -18'd20413;
assign mem3_i[170] = 18'd62276;
assign mem3_r[171] = -18'd18796;
assign mem3_i[171] = 18'd62783;
assign mem3_r[172] = -18'd17166;
assign mem3_i[172] = 18'd63248;
assign mem3_r[173] = -18'd15526;
assign mem3_i[173] = 18'd63670;
assign mem3_r[174] = -18'd13874;
assign mem3_i[174] = 18'd64051;
assign mem3_r[175] = -18'd12214;
assign mem3_i[175] = 18'd64388;
assign mem3_r[176] = -18'd10545;
assign mem3_i[176] = 18'd64682;
assign mem3_r[177] = -18'd8869;
assign mem3_i[177] = 18'd64933;
assign mem3_r[178] = -18'd7187;
assign mem3_i[178] = 18'd65141;
assign mem3_r[179] = -18'd5501;
assign mem3_i[179] = 18'd65305;
assign mem3_r[180] = -18'd3811;
assign mem3_i[180] = 18'd65425;
assign mem3_r[181] = -18'd2118;
assign mem3_i[181] = 18'd65502;
assign mem3_r[182] = -18'd424;
assign mem3_i[182] = 18'd65535;
assign mem3_r[183] = 18'd1271;
assign mem3_i[183] = 18'd65524;
assign mem3_r[184] = 18'd2964;
assign mem3_i[184] = 18'd65469;
assign mem3_r[185] = 18'd4656;
assign mem3_i[185] = 18'd65370;
assign mem3_r[186] = 18'd6345;
assign mem3_i[186] = 18'd65228;
assign mem3_r[187] = 18'd8029;
assign mem3_i[187] = 18'd65042;
assign mem3_r[188] = 18'd9708;
assign mem3_i[188] = 18'd64813;
assign mem3_r[189] = 18'd11380;
assign mem3_i[189] = 18'd64540;
assign mem3_r[190] = 18'd13045;
assign mem3_i[190] = 18'd64225;
assign mem3_r[191] = 18'd14701;
assign mem3_i[191] = 18'd63866;
assign mem3_r[192] = 18'd16347;
assign mem3_i[192] = 18'd63464;
assign mem3_r[193] = 18'd17983;
assign mem3_i[193] = 18'd63021;
assign mem3_r[194] = 18'd19606;
assign mem3_i[194] = 18'd62535;
assign mem3_r[195] = 18'd21216;
assign mem3_i[195] = 18'd62007;
assign mem3_r[196] = 18'd22812;
assign mem3_i[196] = 18'd61438;
assign mem3_r[197] = 18'd24393;
assign mem3_i[197] = 18'd60827;
assign mem3_r[198] = 18'd25957;
assign mem3_i[198] = 18'd60176;
assign mem3_r[199] = 18'd27505;
assign mem3_i[199] = 18'd59485;
assign mem3_r[200] = 18'd29033;
assign mem3_i[200] = 18'd58754;
assign mem3_r[201] = 18'd30543;
assign mem3_i[201] = 18'd57984;
assign mem3_r[202] = 18'd32032;
assign mem3_i[202] = 18'd57175;
assign mem3_r[203] = 18'd33499;
assign mem3_i[203] = 18'd56327;
assign mem3_r[204] = 18'd34944;
assign mem3_i[204] = 18'd55443;
assign mem3_r[205] = 18'd36366;
assign mem3_i[205] = 18'd54521;
assign mem3_r[206] = 18'd37763;
assign mem3_i[206] = 18'd53562;
assign mem3_r[207] = 18'd39135;
assign mem3_i[207] = 18'd52568;
assign mem3_r[208] = 18'd40481;
assign mem3_i[208] = 18'd51539;
assign mem3_r[209] = 18'd41800;
assign mem3_i[209] = 18'd50475;
assign mem3_r[210] = 18'd43091;
assign mem3_i[210] = 18'd49377;
assign mem3_r[211] = 18'd44354;
assign mem3_i[211] = 18'd48247;
assign mem3_r[212] = 18'd45586;
assign mem3_i[212] = 18'd47084;
assign mem3_r[213] = 18'd46788;
assign mem3_i[213] = 18'd45889;
assign mem3_r[214] = 18'd47959;
assign mem3_i[214] = 18'd44664;
assign mem3_r[215] = 18'd49098;
assign mem3_i[215] = 18'd43410;
assign mem3_r[216] = 18'd50203;
assign mem3_i[216] = 18'd42126;
assign mem3_r[217] = 18'd51276;
assign mem3_i[217] = 18'd40814;
assign mem3_r[218] = 18'd52314;
assign mem3_i[218] = 18'd39474;
assign mem3_r[219] = 18'd53317;
assign mem3_i[219] = 18'd38109;
assign mem3_r[220] = 18'd54284;
assign mem3_i[220] = 18'd36717;
assign mem3_r[221] = 18'd55216;
assign mem3_i[221] = 18'd35302;
assign mem3_r[222] = 18'd56110;
assign mem3_i[222] = 18'd33862;
assign mem3_r[223] = 18'd56966;
assign mem3_i[223] = 18'd32400;
assign mem3_r[224] = 18'd57785;
assign mem3_i[224] = 18'd30917;
assign mem3_r[225] = 18'd58565;
assign mem3_i[225] = 18'd29413;
assign mem3_r[226] = 18'd59306;
assign mem3_i[226] = 18'd27889;
assign mem3_r[227] = 18'd60007;
assign mem3_i[227] = 18'd26346;
assign mem3_r[228] = 18'd60668;
assign mem3_i[228] = 18'd24786;
assign mem3_r[229] = 18'd61289;
assign mem3_i[229] = 18'd23209;
assign mem3_r[230] = 18'd61868;
assign mem3_i[230] = 18'd21617;
assign mem3_r[231] = 18'd62407;
assign mem3_i[231] = 18'd20010;
assign mem3_r[232] = 18'd62903;
assign mem3_i[232] = 18'd18390;
assign mem3_r[233] = 18'd63357;
assign mem3_i[233] = 18'd16757;
assign mem3_r[234] = 18'd63769;
assign mem3_i[234] = 18'd15114;
assign mem3_r[235] = 18'd64139;
assign mem3_i[235] = 18'd13460;
assign mem3_r[236] = 18'd64465;
assign mem3_i[236] = 18'd11797;
assign mem3_r[237] = 18'd64749;
assign mem3_i[237] = 18'd10127;
assign mem3_r[238] = 18'd64989;
assign mem3_i[238] = 18'd8449;
assign mem3_r[239] = 18'd65186;
assign mem3_i[239] = 18'd6766;
assign mem3_r[240] = 18'd65339;
assign mem3_i[240] = 18'd5079;
assign mem3_r[241] = 18'd65448;
assign mem3_i[241] = 18'd3388;
assign mem3_r[242] = 18'd65514;
assign mem3_i[242] = 18'd1694;



assign mem2_r[0] = 18'd65536;
assign mem2_i[0] = 18'd0;
assign mem2_r[1] = 18'd65516;
assign mem2_i[1] = -18'd1608;
assign mem2_r[2] = 18'd65457;
assign mem2_i[2] = -18'd3216;
assign mem2_r[3] = 18'd65358;
assign mem2_i[3] = -18'd4821;
assign mem2_r[4] = 18'd65220;
assign mem2_i[4] = -18'd6424;
assign mem2_r[5] = 18'd65043;
assign mem2_i[5] = -18'd8022;
assign mem2_r[6] = 18'd64827;
assign mem2_i[6] = -18'd9616;
assign mem2_r[7] = 18'd64571;
assign mem2_i[7] = -18'd11204;
assign mem2_r[8] = 18'd64277;
assign mem2_i[8] = -18'd12785;
assign mem2_r[9] = 18'd63944;
assign mem2_i[9] = -18'd14359;
assign mem2_r[10] = 18'd63572;
assign mem2_i[10] = -18'd15924;
assign mem2_r[11] = 18'd63162;
assign mem2_i[11] = -18'd17479;
assign mem2_r[12] = 18'd62714;
assign mem2_i[12] = -18'd19024;
assign mem2_r[13] = 18'd62228;
assign mem2_i[13] = -18'd20557;
assign mem2_r[14] = 18'd61705;
assign mem2_i[14] = -18'd22078;
assign mem2_r[15] = 18'd61145;
assign mem2_i[15] = -18'd23586;
assign mem2_r[16] = 18'd60547;
assign mem2_i[16] = -18'd25080;
assign mem2_r[17] = 18'd59914;
assign mem2_i[17] = -18'd26558;
assign mem2_r[18] = 18'd59244;
assign mem2_i[18] = -18'd28020;
assign mem2_r[19] = 18'd58538;
assign mem2_i[19] = -18'd29466;
assign mem2_r[20] = 18'd57798;
assign mem2_i[20] = -18'd30893;
assign mem2_r[21] = 18'd57022;
assign mem2_i[21] = -18'd32303;
assign mem2_r[22] = 18'd56212;
assign mem2_i[22] = -18'd33692;
assign mem2_r[23] = 18'd55368;
assign mem2_i[23] = -18'd35062;
assign mem2_r[24] = 18'd54491;
assign mem2_i[24] = -18'd36410;
assign mem2_r[25] = 18'd53581;
assign mem2_i[25] = -18'd37736;
assign mem2_r[26] = 18'd52639;
assign mem2_i[26] = -18'd39040;
assign mem2_r[27] = 18'd51665;
assign mem2_i[27] = -18'd40320;
assign mem2_r[28] = 18'd50660;
assign mem2_i[28] = -18'd41576;
assign mem2_r[29] = 18'd49624;
assign mem2_i[29] = -18'd42806;
assign mem2_r[30] = 18'd48559;
assign mem2_i[30] = -18'd44011;
assign mem2_r[31] = 18'd47464;
assign mem2_i[31] = -18'd45190;
assign mem2_r[32] = 18'd46341;
assign mem2_i[32] = -18'd46341;
assign mem2_r[33] = 18'd45190;
assign mem2_i[33] = -18'd47464;
assign mem2_r[34] = 18'd44011;
assign mem2_i[34] = -18'd48559;
assign mem2_r[35] = 18'd42806;
assign mem2_i[35] = -18'd49624;
assign mem2_r[36] = 18'd41576;
assign mem2_i[36] = -18'd50660;
assign mem2_r[37] = 18'd40320;
assign mem2_i[37] = -18'd51665;
assign mem2_r[38] = 18'd39040;
assign mem2_i[38] = -18'd52639;
assign mem2_r[39] = 18'd37736;
assign mem2_i[39] = -18'd53581;
assign mem2_r[40] = 18'd36410;
assign mem2_i[40] = -18'd54491;
assign mem2_r[41] = 18'd35062;
assign mem2_i[41] = -18'd55368;
assign mem2_r[42] = 18'd33692;
assign mem2_i[42] = -18'd56212;
assign mem2_r[43] = 18'd32303;
assign mem2_i[43] = -18'd57022;
assign mem2_r[44] = 18'd30893;
assign mem2_i[44] = -18'd57798;
assign mem2_r[45] = 18'd29466;
assign mem2_i[45] = -18'd58538;
assign mem2_r[46] = 18'd28020;
assign mem2_i[46] = -18'd59244;
assign mem2_r[47] = 18'd26558;
assign mem2_i[47] = -18'd59914;
assign mem2_r[48] = 18'd25080;
assign mem2_i[48] = -18'd60547;
assign mem2_r[49] = 18'd23586;
assign mem2_i[49] = -18'd61145;
assign mem2_r[50] = 18'd22078;
assign mem2_i[50] = -18'd61705;
assign mem2_r[51] = 18'd20557;
assign mem2_i[51] = -18'd62228;
assign mem2_r[52] = 18'd19024;
assign mem2_i[52] = -18'd62714;
assign mem2_r[53] = 18'd17479;
assign mem2_i[53] = -18'd63162;
assign mem2_r[54] = 18'd15924;
assign mem2_i[54] = -18'd63572;
assign mem2_r[55] = 18'd14359;
assign mem2_i[55] = -18'd63944;
assign mem2_r[56] = 18'd12785;
assign mem2_i[56] = -18'd64277;
assign mem2_r[57] = 18'd11204;
assign mem2_i[57] = -18'd64571;
assign mem2_r[58] = 18'd9616;
assign mem2_i[58] = -18'd64827;
assign mem2_r[59] = 18'd8022;
assign mem2_i[59] = -18'd65043;
assign mem2_r[60] = 18'd6424;
assign mem2_i[60] = -18'd65220;
assign mem2_r[61] = 18'd4821;
assign mem2_i[61] = -18'd65358;
assign mem2_r[62] = 18'd3216;
assign mem2_i[62] = -18'd65457;
assign mem2_r[63] = 18'd1608;
assign mem2_i[63] = -18'd65516;
assign mem2_r[64] = 18'd0;
assign mem2_i[64] = -18'd65536;
assign mem2_r[65] = -18'd1608;
assign mem2_i[65] = -18'd65516;
assign mem2_r[66] = -18'd3216;
assign mem2_i[66] = -18'd65457;
assign mem2_r[67] = -18'd4821;
assign mem2_i[67] = -18'd65358;
assign mem2_r[68] = -18'd6424;
assign mem2_i[68] = -18'd65220;
assign mem2_r[69] = -18'd8022;
assign mem2_i[69] = -18'd65043;
assign mem2_r[70] = -18'd9616;
assign mem2_i[70] = -18'd64827;
assign mem2_r[71] = -18'd11204;
assign mem2_i[71] = -18'd64571;
assign mem2_r[72] = -18'd12785;
assign mem2_i[72] = -18'd64277;
assign mem2_r[73] = -18'd14359;
assign mem2_i[73] = -18'd63944;
assign mem2_r[74] = -18'd15924;
assign mem2_i[74] = -18'd63572;
assign mem2_r[75] = -18'd17479;
assign mem2_i[75] = -18'd63162;
assign mem2_r[76] = -18'd19024;
assign mem2_i[76] = -18'd62714;
assign mem2_r[77] = -18'd20557;
assign mem2_i[77] = -18'd62228;
assign mem2_r[78] = -18'd22078;
assign mem2_i[78] = -18'd61705;
assign mem2_r[79] = -18'd23586;
assign mem2_i[79] = -18'd61145;
assign mem2_r[80] = -18'd25080;
assign mem2_i[80] = -18'd60547;
assign mem2_r[81] = -18'd26558;
assign mem2_i[81] = -18'd59914;
assign mem2_r[82] = -18'd28020;
assign mem2_i[82] = -18'd59244;
assign mem2_r[83] = -18'd29466;
assign mem2_i[83] = -18'd58538;
assign mem2_r[84] = -18'd30893;
assign mem2_i[84] = -18'd57798;
assign mem2_r[85] = -18'd32303;
assign mem2_i[85] = -18'd57022;
assign mem2_r[86] = -18'd33692;
assign mem2_i[86] = -18'd56212;
assign mem2_r[87] = -18'd35062;
assign mem2_i[87] = -18'd55368;
assign mem2_r[88] = -18'd36410;
assign mem2_i[88] = -18'd54491;
assign mem2_r[89] = -18'd37736;
assign mem2_i[89] = -18'd53581;
assign mem2_r[90] = -18'd39040;
assign mem2_i[90] = -18'd52639;
assign mem2_r[91] = -18'd40320;
assign mem2_i[91] = -18'd51665;
assign mem2_r[92] = -18'd41576;
assign mem2_i[92] = -18'd50660;
assign mem2_r[93] = -18'd42806;
assign mem2_i[93] = -18'd49624;
assign mem2_r[94] = -18'd44011;
assign mem2_i[94] = -18'd48559;
assign mem2_r[95] = -18'd45190;
assign mem2_i[95] = -18'd47464;
assign mem2_r[96] = -18'd46341;
assign mem2_i[96] = -18'd46341;
assign mem2_r[97] = -18'd47464;
assign mem2_i[97] = -18'd45190;
assign mem2_r[98] = -18'd48559;
assign mem2_i[98] = -18'd44011;
assign mem2_r[99] = -18'd49624;
assign mem2_i[99] = -18'd42806;
assign mem2_r[100] = -18'd50660;
assign mem2_i[100] = -18'd41576;
assign mem2_r[101] = -18'd51665;
assign mem2_i[101] = -18'd40320;
assign mem2_r[102] = -18'd52639;
assign mem2_i[102] = -18'd39040;
assign mem2_r[103] = -18'd53581;
assign mem2_i[103] = -18'd37736;
assign mem2_r[104] = -18'd54491;
assign mem2_i[104] = -18'd36410;
assign mem2_r[105] = -18'd55368;
assign mem2_i[105] = -18'd35062;
assign mem2_r[106] = -18'd56212;
assign mem2_i[106] = -18'd33692;
assign mem2_r[107] = -18'd57022;
assign mem2_i[107] = -18'd32303;
assign mem2_r[108] = -18'd57798;
assign mem2_i[108] = -18'd30893;
assign mem2_r[109] = -18'd58538;
assign mem2_i[109] = -18'd29466;
assign mem2_r[110] = -18'd59244;
assign mem2_i[110] = -18'd28020;
assign mem2_r[111] = -18'd59914;
assign mem2_i[111] = -18'd26558;
assign mem2_r[112] = -18'd60547;
assign mem2_i[112] = -18'd25080;
assign mem2_r[113] = -18'd61145;
assign mem2_i[113] = -18'd23586;
assign mem2_r[114] = -18'd61705;
assign mem2_i[114] = -18'd22078;
assign mem2_r[115] = -18'd62228;
assign mem2_i[115] = -18'd20557;
assign mem2_r[116] = -18'd62714;
assign mem2_i[116] = -18'd19024;
assign mem2_r[117] = -18'd63162;
assign mem2_i[117] = -18'd17479;
assign mem2_r[118] = -18'd63572;
assign mem2_i[118] = -18'd15924;
assign mem2_r[119] = -18'd63944;
assign mem2_i[119] = -18'd14359;
assign mem2_r[120] = -18'd64277;
assign mem2_i[120] = -18'd12785;
assign mem2_r[121] = -18'd64571;
assign mem2_i[121] = -18'd11204;
assign mem2_r[122] = -18'd64827;
assign mem2_i[122] = -18'd9616;
assign mem2_r[123] = -18'd65043;
assign mem2_i[123] = -18'd8022;
assign mem2_r[124] = -18'd65220;
assign mem2_i[124] = -18'd6424;
assign mem2_r[125] = -18'd65358;
assign mem2_i[125] = -18'd4821;
assign mem2_r[126] = -18'd65457;
assign mem2_i[126] = -18'd3216;
assign mem2_r[127] = -18'd65516;
assign mem2_i[127] = -18'd1608;
assign mem2_r[128] = -18'd65536;
assign mem2_i[128] = 18'd0;
assign mem2_r[129] = -18'd65516;
assign mem2_i[129] = 18'd1608;
assign mem2_r[130] = -18'd65457;
assign mem2_i[130] = 18'd3216;
assign mem2_r[131] = -18'd65358;
assign mem2_i[131] = 18'd4821;
assign mem2_r[132] = -18'd65220;
assign mem2_i[132] = 18'd6424;
assign mem2_r[133] = -18'd65043;
assign mem2_i[133] = 18'd8022;
assign mem2_r[134] = -18'd64827;
assign mem2_i[134] = 18'd9616;
assign mem2_r[135] = -18'd64571;
assign mem2_i[135] = 18'd11204;
assign mem2_r[136] = -18'd64277;
assign mem2_i[136] = 18'd12785;
assign mem2_r[137] = -18'd63944;
assign mem2_i[137] = 18'd14359;
assign mem2_r[138] = -18'd63572;
assign mem2_i[138] = 18'd15924;
assign mem2_r[139] = -18'd63162;
assign mem2_i[139] = 18'd17479;
assign mem2_r[140] = -18'd62714;
assign mem2_i[140] = 18'd19024;
assign mem2_r[141] = -18'd62228;
assign mem2_i[141] = 18'd20557;
assign mem2_r[142] = -18'd61705;
assign mem2_i[142] = 18'd22078;
assign mem2_r[143] = -18'd61145;
assign mem2_i[143] = 18'd23586;
assign mem2_r[144] = -18'd60547;
assign mem2_i[144] = 18'd25080;
assign mem2_r[145] = -18'd59914;
assign mem2_i[145] = 18'd26558;
assign mem2_r[146] = -18'd59244;
assign mem2_i[146] = 18'd28020;
assign mem2_r[147] = -18'd58538;
assign mem2_i[147] = 18'd29466;
assign mem2_r[148] = -18'd57798;
assign mem2_i[148] = 18'd30893;
assign mem2_r[149] = -18'd57022;
assign mem2_i[149] = 18'd32303;
assign mem2_r[150] = -18'd56212;
assign mem2_i[150] = 18'd33692;
assign mem2_r[151] = -18'd55368;
assign mem2_i[151] = 18'd35062;
assign mem2_r[152] = -18'd54491;
assign mem2_i[152] = 18'd36410;
assign mem2_r[153] = -18'd53581;
assign mem2_i[153] = 18'd37736;
assign mem2_r[154] = -18'd52639;
assign mem2_i[154] = 18'd39040;
assign mem2_r[155] = -18'd51665;
assign mem2_i[155] = 18'd40320;
assign mem2_r[156] = -18'd50660;
assign mem2_i[156] = 18'd41576;
assign mem2_r[157] = -18'd49624;
assign mem2_i[157] = 18'd42806;
assign mem2_r[158] = -18'd48559;
assign mem2_i[158] = 18'd44011;
assign mem2_r[159] = -18'd47464;
assign mem2_i[159] = 18'd45190;
assign mem2_r[160] = -18'd46341;
assign mem2_i[160] = 18'd46341;
assign mem2_r[161] = -18'd45190;
assign mem2_i[161] = 18'd47464;
assign mem2_r[162] = -18'd44011;
assign mem2_i[162] = 18'd48559;
assign mem2_r[163] = -18'd42806;
assign mem2_i[163] = 18'd49624;
assign mem2_r[164] = -18'd41576;
assign mem2_i[164] = 18'd50660;
assign mem2_r[165] = -18'd40320;
assign mem2_i[165] = 18'd51665;
assign mem2_r[166] = -18'd39040;
assign mem2_i[166] = 18'd52639;
assign mem2_r[167] = -18'd37736;
assign mem2_i[167] = 18'd53581;
assign mem2_r[168] = -18'd36410;
assign mem2_i[168] = 18'd54491;
assign mem2_r[169] = -18'd35062;
assign mem2_i[169] = 18'd55368;
assign mem2_r[170] = -18'd33692;
assign mem2_i[170] = 18'd56212;
assign mem2_r[171] = -18'd32303;
assign mem2_i[171] = 18'd57022;
assign mem2_r[172] = -18'd30893;
assign mem2_i[172] = 18'd57798;
assign mem2_r[173] = -18'd29466;
assign mem2_i[173] = 18'd58538;
assign mem2_r[174] = -18'd28020;
assign mem2_i[174] = 18'd59244;
assign mem2_r[175] = -18'd26558;
assign mem2_i[175] = 18'd59914;
assign mem2_r[176] = -18'd25080;
assign mem2_i[176] = 18'd60547;
assign mem2_r[177] = -18'd23586;
assign mem2_i[177] = 18'd61145;
assign mem2_r[178] = -18'd22078;
assign mem2_i[178] = 18'd61705;
assign mem2_r[179] = -18'd20557;
assign mem2_i[179] = 18'd62228;
assign mem2_r[180] = -18'd19024;
assign mem2_i[180] = 18'd62714;
assign mem2_r[181] = -18'd17479;
assign mem2_i[181] = 18'd63162;
assign mem2_r[182] = -18'd15924;
assign mem2_i[182] = 18'd63572;
assign mem2_r[183] = -18'd14359;
assign mem2_i[183] = 18'd63944;
assign mem2_r[184] = -18'd12785;
assign mem2_i[184] = 18'd64277;
assign mem2_r[185] = -18'd11204;
assign mem2_i[185] = 18'd64571;
assign mem2_r[186] = -18'd9616;
assign mem2_i[186] = 18'd64827;
assign mem2_r[187] = -18'd8022;
assign mem2_i[187] = 18'd65043;
assign mem2_r[188] = -18'd6424;
assign mem2_i[188] = 18'd65220;
assign mem2_r[189] = -18'd4821;
assign mem2_i[189] = 18'd65358;
assign mem2_r[190] = -18'd3216;
assign mem2_i[190] = 18'd65457;
assign mem2_r[191] = -18'd1608;
assign mem2_i[191] = 18'd65516;
assign mem2_r[192] = 18'd0;
assign mem2_i[192] = 18'd65536;
assign mem2_r[193] = 18'd1608;
assign mem2_i[193] = 18'd65516;
assign mem2_r[194] = 18'd3216;
assign mem2_i[194] = 18'd65457;
assign mem2_r[195] = 18'd4821;
assign mem2_i[195] = 18'd65358;
assign mem2_r[196] = 18'd6424;
assign mem2_i[196] = 18'd65220;
assign mem2_r[197] = 18'd8022;
assign mem2_i[197] = 18'd65043;
assign mem2_r[198] = 18'd9616;
assign mem2_i[198] = 18'd64827;
assign mem2_r[199] = 18'd11204;
assign mem2_i[199] = 18'd64571;
assign mem2_r[200] = 18'd12785;
assign mem2_i[200] = 18'd64277;
assign mem2_r[201] = 18'd14359;
assign mem2_i[201] = 18'd63944;
assign mem2_r[202] = 18'd15924;
assign mem2_i[202] = 18'd63572;
assign mem2_r[203] = 18'd17479;
assign mem2_i[203] = 18'd63162;
assign mem2_r[204] = 18'd19024;
assign mem2_i[204] = 18'd62714;
assign mem2_r[205] = 18'd20557;
assign mem2_i[205] = 18'd62228;
assign mem2_r[206] = 18'd22078;
assign mem2_i[206] = 18'd61705;
assign mem2_r[207] = 18'd23586;
assign mem2_i[207] = 18'd61145;
assign mem2_r[208] = 18'd25080;
assign mem2_i[208] = 18'd60547;
assign mem2_r[209] = 18'd26558;
assign mem2_i[209] = 18'd59914;
assign mem2_r[210] = 18'd28020;
assign mem2_i[210] = 18'd59244;
assign mem2_r[211] = 18'd29466;
assign mem2_i[211] = 18'd58538;
assign mem2_r[212] = 18'd30893;
assign mem2_i[212] = 18'd57798;
assign mem2_r[213] = 18'd32303;
assign mem2_i[213] = 18'd57022;
assign mem2_r[214] = 18'd33692;
assign mem2_i[214] = 18'd56212;
assign mem2_r[215] = 18'd35062;
assign mem2_i[215] = 18'd55368;
assign mem2_r[216] = 18'd36410;
assign mem2_i[216] = 18'd54491;
assign mem2_r[217] = 18'd37736;
assign mem2_i[217] = 18'd53581;
assign mem2_r[218] = 18'd39040;
assign mem2_i[218] = 18'd52639;
assign mem2_r[219] = 18'd40320;
assign mem2_i[219] = 18'd51665;
assign mem2_r[220] = 18'd41576;
assign mem2_i[220] = 18'd50660;
assign mem2_r[221] = 18'd42806;
assign mem2_i[221] = 18'd49624;
assign mem2_r[222] = 18'd44011;
assign mem2_i[222] = 18'd48559;
assign mem2_r[223] = 18'd45190;
assign mem2_i[223] = 18'd47464;
assign mem2_r[224] = 18'd46341;
assign mem2_i[224] = 18'd46341;
assign mem2_r[225] = 18'd47464;
assign mem2_i[225] = 18'd45190;
assign mem2_r[226] = 18'd48559;
assign mem2_i[226] = 18'd44011;
assign mem2_r[227] = 18'd49624;
assign mem2_i[227] = 18'd42806;
assign mem2_r[228] = 18'd50660;
assign mem2_i[228] = 18'd41576;
assign mem2_r[229] = 18'd51665;
assign mem2_i[229] = 18'd40320;
assign mem2_r[230] = 18'd52639;
assign mem2_i[230] = 18'd39040;
assign mem2_r[231] = 18'd53581;
assign mem2_i[231] = 18'd37736;
assign mem2_r[232] = 18'd54491;
assign mem2_i[232] = 18'd36410;
assign mem2_r[233] = 18'd55368;
assign mem2_i[233] = 18'd35062;
assign mem2_r[234] = 18'd56212;
assign mem2_i[234] = 18'd33692;
assign mem2_r[235] = 18'd57022;
assign mem2_i[235] = 18'd32303;
assign mem2_r[236] = 18'd57798;
assign mem2_i[236] = 18'd30893;
assign mem2_r[237] = 18'd58538;
assign mem2_i[237] = 18'd29466;
assign mem2_r[238] = 18'd59244;
assign mem2_i[238] = 18'd28020;
assign mem2_r[239] = 18'd59914;
assign mem2_i[239] = 18'd26558;
assign mem2_r[240] = 18'd60547;
assign mem2_i[240] = 18'd25080;
assign mem2_r[241] = 18'd61145;
assign mem2_i[241] = 18'd23586;
assign mem2_r[242] = 18'd61705;
assign mem2_i[242] = 18'd22078;
assign mem2_r[243] = 18'd62228;
assign mem2_i[243] = 18'd20557;
assign mem2_r[244] = 18'd62714;
assign mem2_i[244] = 18'd19024;
assign mem2_r[245] = 18'd63162;
assign mem2_i[245] = 18'd17479;
assign mem2_r[246] = 18'd63572;
assign mem2_i[246] = 18'd15924;
assign mem2_r[247] = 18'd63944;
assign mem2_i[247] = 18'd14359;
assign mem2_r[248] = 18'd64277;
assign mem2_i[248] = 18'd12785;
assign mem2_r[249] = 18'd64571;
assign mem2_i[249] = 18'd11204;
assign mem2_r[250] = 18'd64827;
assign mem2_i[250] = 18'd9616;
assign mem2_r[251] = 18'd65043;
assign mem2_i[251] = 18'd8022;
assign mem2_r[252] = 18'd65220;
assign mem2_i[252] = 18'd6424;
assign mem2_r[253] = 18'd65358;
assign mem2_i[253] = 18'd4821;
assign mem2_r[254] = 18'd65457;
assign mem2_i[254] = 18'd3216;
assign mem2_r[255] = 18'd65516;
assign mem2_i[255] = 18'd1608;




endmodule